//////////////////////////////////////////////////////////////////////////////
// hw2_prob1.sv
//
// Author:	Alex Beaulier (roy.kravitz@pdx.edu)
// Date:	9-5-2020 (modified 9-5-2021)
//
// Contains instantiation of top level model ALU and includes register file. 
// 
/////////////////////////////////////////////////////////////////////////////
